parameter string g_data_dir_path = "/work/kam/srup_dpi_core_test/data";
